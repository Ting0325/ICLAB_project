module reorder_buff(
	input inst
	
);



endmodule
