/*
 * keeps track of which reservation station a register is waiting on
 *
 *
 * */

module rename_tbl(

);

endmodule
